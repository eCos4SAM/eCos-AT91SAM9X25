# ====================================================================
#
#      hal_arm_at91_sam7s.cdl
#
#      ARM AT91 SAM7 HAL package configuration data
#
# ====================================================================
## ####ECOSGPLCOPYRIGHTBEGIN####                                            
## -------------------------------------------                              
## This file is part of eCos, the Embedded Configurable Operating System.   
## Copyright (C) 1998, 1999, 2000, 2001, 2002, 2003, 2005 Free Software Foundation, Inc.
##
## eCos is free software; you can redistribute it and/or modify it under    
## the terms of the GNU General Public License as published by the Free     
## Software Foundation; either version 2 or (at your option) any later      
## version.                                                                 
##
## eCos is distributed in the hope that it will be useful, but WITHOUT      
## ANY WARRANTY; without even the implied warranty of MERCHANTABILITY or    
## FITNESS FOR A PARTICULAR PURPOSE.  See the GNU General Public License    
## for more details.                                                        
##
## You should have received a copy of the GNU General Public License        
## along with eCos; if not, write to the Free Software Foundation, Inc.,    
## 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.            
##
## As a special exception, if other files instantiate templates or use      
## macros or inline functions from this file, or you compile this file      
## and link it with other works to produce a work based on this file,       
## this file does not by itself cause the resulting work to be covered by   
## the GNU General Public License. However the source code for this file    
## must still be made available in accordance with section (3) of the GNU   
## General Public License v2.                                               
##
## This exception does not invalidate any other reasons why a work based    
## on this file might be covered by the GNU General Public License.         
## -------------------------------------------                              
## ####ECOSGPLCOPYRIGHTEND####                                              
# ====================================================================
######DESCRIPTIONBEGIN####
#
# Author(s):      Owen Kirby
# Contributors:   
# Date:           2009-11-12
#
#####DESCRIPTIONEND####
#
# ====================================================================

# =============================================================================
# Key-change    Date       Author   Description
# --------------+----------+--------+------------------------------------------
# SAM9X25-0001  2011/03/20 TuPN     Create new platform sam9x25 (base on g20)
# SAM9G45-0001  2011/03/20 TuPN     Create new platform sam9g45 (base on g20)
#
#==============================================================================

cdl_package CYGPKG_HAL_ARM_AT91SAM9 {
    display       "Atmel AT91SAM9 HAL"
    parent        CYGPKG_HAL_ARM
    define_header hal_arm_at91sam9.h
    include_dir   cyg/hal
    hardware
    description   "
        The AT91SAM9 HAL package provides the support needed to run
        eCos on an Atmel AT91SAM9 based board."

    compile       at91sam9_misc.c
    
    requires      { CYGHWR_HAL_ARM_AT91_FIQ     }

    implements    CYGINT_HAL_ARM_AT91_SERIAL_DBG_HW
    implements    CYGINT_HAL_ARM_AT91_PIT_HW
    implements    CYGINT_HAL_ARM_AT91_SYS_INTERRUPT

    define_proc {
        puts $::cdl_system_header "#define CYGBLD_HAL_TARGET_H   <pkgconf/hal_arm.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_VARIANT_H  <pkgconf/hal_arm_at91.h>"
        puts $::cdl_system_header "#define CYGBLD_HAL_ARM_VAR_IO_H"
    }

    cdl_option CYGHWR_HAL_ARM_AT91SAM9 {
        display        "AT91SAM9 variant used"
        flavor         data
        default_value  {"at91sam9g20"}
#SAM9X25-0001.DEL        legal_values   {"at91sam9g10" "at91sam9g20" "at91sam9g45" }
#SAM9X25-0001.ADD.Start
#SAM9G45-0001.Modified.Start
        legal_values   {"at91sam9g10" "at91sam9g20"
                 		"at91sam9g45"
						"at91sam9x25"	}
#SAM9G45-0001.Modified.End
#SAM9X25-0001.ADD.End
        description    "
           The AT91SAM9 microcontroller family has several variants,
           the main differences being the amount of on-chip SRAM,
           FLASH, peripherals and their layout. This option allows the
           platform HALs to select the specific microcontroller
           being used."
    }

    cdl_option CYGBLD_HAL_ARM_AT91SAM9_USB {
        display       "USB device"
#SAM9X25-0001.DEL        active_if     { CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g10" ||
#SAM9X25-0001.DEL                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g20" ||
#SAM9X25-0001.DEL                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g45" }
#SAM9X25-0001.ADD.Start
        active_if     { CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g10" ||
                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g20" ||
                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g45" ||
                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9x25" 
                      }
#SAM9X25-0001.ADD.End                        
                                                
        implements    CYGINT_DEVS_USB_AT91_HAS_USB
        default_value 1
        no_define
        description   "
            All but the AT91SAM7S32 has the USB device"
    }

    cdl_option CYGBLD_HAL_ARM_AT91SAM9_SPI1 {
        display       "Second SPI bus controller"
#SAM9X25-0001.DEL        active_if     { CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g10" ||
#SAM9X25-0001.DEL                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g20" ||
#SAM9X25-0001.DEL                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g45" }
#SAM9X25-0001.ADD.Start
        active_if     { CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g10" ||
                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g20" ||
                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9g45" ||
                        CYGHWR_HAL_ARM_AT91SAM9 == "at91sam9x25"
                      }
#SAM9X25-0001.ADD.End
                        
        implements    CYGINT_DEVS_SPI_ARM_AT91_HAS_BUS1
        default_value 1
        no_define
        description   "
            The SAM7X and SAM7XC have the second SPI bus controller"
    }

    cdl_component CYGNUM_HAL_RTC_CONSTANTS {
        display       "Real-time clock constants"
        flavor        none

        cdl_option CYGNUM_HAL_RTC_NUMERATOR {
            display       "Real-time clock numerator"
            flavor        data
            default_value 1000000000
        }
        cdl_option CYGNUM_HAL_RTC_DENOMINATOR {
            display       "Real-time clock denominator"
            flavor        data
            default_value 100
        }
        cdl_option CYGNUM_HAL_RTC_PERIOD {
            display       "Real-time clock period"
            flavor        data
#SAM9X25-0001.DEL legal_values  1 to 0xffff
#SAM9X25-0001.ADD.Start
			legal_values  1 to (CYGBLD_HAL_ARM_AT91_TIMER_TC ? 0xffff : 0xfffff)
#SAM9X25-0001.ADD.End
            calculated    { (CYGNUM_HAL_RTC_NUMERATOR * 
                             CYGNUM_HAL_ARM_AT91_CLOCK_SPEED /
                             (CYGBLD_HAL_ARM_AT91_TIMER_TC ? 32 : 16) / 
                             CYGNUM_HAL_RTC_DENOMINATOR / 
                             1000000000
                            )
                          }
            description   "Value to program into the RTC clock generator."
        }
    }
    
    cdl_component CYG_HAL_STARTUP {
        display       "Startup type"
        flavor        data
        default_value {"RAM"}
        legal_values  {"RAM"}
        no_define
        define -file system.h CYG_HAL_STARTUP
        description   "
            When targeting the AT91SAM9 eval boards it is possible to build
            the system for either RAM bootstrap or ROM bootstrap(s). Select
            'ram' when building programs to load into RAM using on board
            debug software such as Angel or eCos GDB stubs.  Select 'rom'
            when building a stand-alone application which will be put
            into ROM"
    }

    # Real-time clock/counter specifics
    cdl_option CYGNUM_HAL_ARM_AT91_CLOCK_SPEED {
        display       "CPU clock speed"
        flavor        data
        calculated    { CYGNUM_HAL_ARM_AT91_CLOCK_OSC_MAIN *
                        CYGNUM_HAL_ARM_AT91_PLL_MULTIPLIER /
                        CYGNUM_HAL_ARM_AT91_PLL_DIVIDER / 2}
        legal_values  { 0 to 220000000 }
        description   "
            The master clock-frequency has to be 48MHz, 96MHz or
            192MHz for the USB to work correctly. The clock setup uses
            PLL clock divided by two"
    }

    cdl_option CYGNUM_HAL_ARM_AT91_CLOCK_XIN_FREQ_MAX {
        display       "Input clock frequency maximum"
        flavor        data
        calculated    { CYGNUM_HAL_ARM_AT91_CLOCK_TYPE == "CRYSTAL" ? 
                        20000000 : 50000000 }
        description   "

            The oscilator in the AT91SAM allows a crystal of up to
            20MHz. However by feeding in directly a clock signal, it
            is possible to use upto 50MHz in XIN."
     }

    cdl_option CYGNUM_HAL_ARM_AT91_CLOCK_OSC_MAIN {
        display       "Main oscillator frequency"
        flavor        data
        legal_values  { 3000000 to CYGNUM_HAL_ARM_AT91_CLOCK_XIN_FREQ_MAX } 
#SAM9X25-0001.ADD.Del default_value { 18432000 }
#SAM9X25-0001.ADD.Start
		default_value { 12000000 }
#SAM9X25-0001.ADD.End
        description   "
            The frequency of the clock input, be it a crystal or a clock 
            signal"
    }

    cdl_option CYGNUM_HAL_ARM_AT91_CLOCK_TYPE {
        display       "Type of main frequency input"
        flavor        data
        default_value { "CRYSTAL" }
        legal_values  { "CRYSTAL" "EXTCLOCK" } 
        description   "
            Whether a crystal or a XIN input clock is clocking the device."
    }

    cdl_option CYGNUM_HAL_ARM_AT91_PMC_MOR_OSCCOUNT {
        display       "Startup time for the main oscillator"
        flavor        data
        legal_values  { 0 to 255 }
        default_value 64
        description   "
            Specifies the number of Slow Clock cycles multiplied by 8 
	    for the Main Oscillator start-up time. 64 is the number suggested
	    by the kind folk at Atmel"
    }       

    cdl_option CYGNUM_HAL_ARM_AT91_PLL_DIVIDER {
        display       "Divider for PLL clock"
        flavor        data
        legal_values  { 0 to 255 }
#SAM9X25-0001.ADD.Del default_value 3
#SAM9X25-0001.ADD.Start
		default_value 9
#SAM9X25-0001.ADD.Start
        description   "
            The X-tal clock is divided by this value when generating the
            PLL clock"
    }       
        
    cdl_option CYGNUM_HAL_ARM_AT91_PLL_MULTIPLIER {
        display       "Multiplier for PLL clock"
        flavor        data
        legal_values  { 0 to 2047 }
#SAM9X25-0001.ADD.Del default_value 43
#SAM9X25-0001.ADD.Start
		default_value 200
#SAM9X25-0001.ADD.Start
        description   "
           The X-tal clock is multiplied by this value when generating
           the PLL clock."
    }

    cdl_option CYGNUM_HAL_ARM_AT91_PLL_COUNT {
        display       "Startup Counter for PLL clock"
        flavor        data
        legal_values  { 0 to 64 }
        default_value 16
        description   "
            Specifies the number of slow clock cycles before the LOCK bit 
	    is set in PMC_SR after PLL Register is written. The Atmel people
	    suggest that 16 should be fine"
    }       
    
    cdl_option CYGNUM_HAL_ARM_AT91_SLOW_CLOCK {
        display       "Slow clock frequency"
        flavor        data
        default_value { 32768 }
        description   "
            The slow clock is an LC oscillator which runs all the
            time. The accuracy of this clock is not very high and 
            is temperature dependent."
    }

    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS {
        display       "Number of communication channels on the board"
        flavor        data
        default_value 3
        description   "
            The AT91SAM9G20-EK has three serial ports, USART0, USART1 and the
            debug port mapped to USART2."
    }
#SAM9X25-0001.TBD.Start
# Need check for x25 & g20
# Need check for g45 & g20
#SAM9X25-0001.TBD.End
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL {
        display          "Debug serial port"
        active_if        CYGPRI_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_CONFIGURABLE
        flavor data
        legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
        default_value    1
        description      "
            The AT91SAM79G20-EK has three serial ports. This option
            chooses which port will be used to connect to a host
            running GDB."
     }
 
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL {
         display          "Diagnostic serial port"
         active_if        CYGPRI_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_CONFIGURABLE
         flavor data
         legal_values     0 to CYGNUM_HAL_VIRTUAL_VECTOR_COMM_CHANNELS-1
         default_value    2
         description      "
            The AT91SAM7S board has three USART serial ports. This option
            chooses which port will be used for diagnostic output."
     }
     
     cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_CONSOLE_CHANNEL_BAUD {
        display       "Diagnostic serial port baud rate"
        flavor        data
        legal_values  9600 19200 38400 57600 115200
        default_value 115200
        description   "
            This option selects the baud rate used for the diagnostic port."
    }
 
    cdl_option CYGNUM_HAL_VIRTUAL_VECTOR_DEBUG_CHANNEL_BAUD {
         display       "GDB serial port baud rate"
         flavor        data
         legal_values  9600 19200 38400 57600 115200
         default_value 38400
         description   "
            This option controls the baud rate used for the GDB connection."
     }
 
    cdl_option CYGBLD_HAL_ARM_AT91_BAUD_DYNAMIC {
        display       "Dynamic calculation of baud rate"
        default_value 0
        description   "
             The AT91SAM7S has a flexible clock generation mechanism 
             where the main clock used to drive peripherals can be
             changed during run time. Such changes affect the serial port
             baud rate generators. Enabling this option includes code 
             which calculates the baud rate setting dynamically from the
             current clock settings. Without this option a static
             calculation is performed which assumes the clock frequency
             has not been changed."
    }

    cdl_component CYGBLD_GLOBAL_OPTIONS {
        display "Global build options"
        flavor  none
        parent  CYGPKG_NONE
        description   "
            Global build options including control over
            compiler flags, linker flags and choice of toolchain."

        cdl_option CYGBLD_GLOBAL_COMMAND_PREFIX {
            display "Global command prefix"
            flavor  data
            no_define
            default_value { "arm-none-eabi" }
            description "
                This option specifies the command prefix used when
                invoking the build tools."
        }

        cdl_option CYGBLD_GLOBAL_CFLAGS {
            display "Global compiler flags"
            flavor  data
            no_define
            default_value { CYGBLD_GLOBAL_WARNFLAGS . CYGBLD_ARCH_CFLAGS .
                            "-mcpu=arm926ej-s -msoft-float -g -O2 -ffunction-sections -fdata-sections -fno-rtti -fno-exceptions -fvtable-gc -finit-priority" }
            description   "
                This option controls the global compiler flags which are used to
                compile all packages by default. Individual packages may define
                options which override these global flags."
        }

        cdl_option CYGBLD_GLOBAL_LDFLAGS {
            display "Global linker flags"
            flavor  data
            no_define
            default_value { CYGBLD_ARCH_LDFLAGS . "-mcpu=arm926ej-s -msoft-float -Wl,--gc-sections -Wl,-static -g -nostdlib" }
            description   "
                This option controls the global linker flags. Individual
                packages may define options which override these global flags."
        }
    }
}
